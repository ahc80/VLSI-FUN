// 

module red (
    
);