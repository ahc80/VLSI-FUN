module speaker ();
    initial begin
        $display("I am speaker!");
    end
endmodule