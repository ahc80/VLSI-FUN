library ieee;
use ieee.std._logic_1164.all;

