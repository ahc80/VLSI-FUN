module txfifo (
    input        PSEL,
    input        PWRITE,
    input        CLEAR_B,
    input        PCLK,
    input  [7:0] TxData,
    output [7:0] PWDATA
);
    
endmodule