module long_divider (
    input[3:0] M,
    input[3:0] D,
    
);
    
endmodule