module proto_tab_tb ();
    
    
endmodule