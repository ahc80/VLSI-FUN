module and_of_gate (
    input  A,
    input  B,
    output S
);

assign S = A & B;
    
endmodule