module ssp (
    ports
);
    
endmodule