module rxfifo (
    input        PSEL,
    input        PWRITE,
    input  [7:0] PWDATA,
    input        CLEAR_B,
    input        PCLK,
    output       SSPTXINTR,
    output [7:0] TxData
);
    
endmodule