module concaternator_dynamic (
    input [1:0]
);
    
endmodule